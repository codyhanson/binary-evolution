/*
Module:			

Description:		

Hierarchy:		


Team Binary Evolution
Ben Fuhrmann, Cody Hanson, Eric Harris, Ross Nordstrom, Eric Weisman

Module designed by:	
Edited by:		
Module interface by:	

Date:			

*/

module template(input clk, 
			  input rst,
			  input
			  output );

	

endmodule;